//module	instructionsBitMap	(	
//			input	logic	clk,
//			input	logic	resetN,
//			input logic	[10:0] offsetX,// offset from top left  position 
//			input logic	[10:0] offsetY,
//			input	logic	InsideRectangle, //input that the pixel is within a bracket 
//)

