// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	StatsDisplayBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,// offset from top left  position 
					input logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic [3:0] level,
					input logic [3:0] birdsLeft,
					input logic [11:0] score,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 

parameter  logic	[7:0] text_color = 8'h00 ; //set the color of the digit 


logic [0:15] [3:0]  MazeBitMapMask ;  

// 8 - level number (based on input)
// 9 - number of birds left (based on input)
// A - level label "L"
// B - level label "v."
// C - heart label
// 3 - score digit (based on input)
// 4 - score digit (based on input)
// 5 - score digit (based on input)
// 6 - score digit (based on input)
logic [0:15] [3:0]  MazeDefaultBitMapMask= 64'hAB80009C0003456000;
 
 
bit [0:9] [0:31] [0:31] number_bitmap  = {
        {
				32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000,
            32'b00000011111111111111111111000000,
            32'b00001111111111111111111111110000,
            32'b00011111111111111111111111111000,
            32'b00111111111111111111111111111100,
            32'b01111111111111111111111111111110,
            32'b11111111111000000000111111111111,
            32'b11111111110000000000011111111111,
            32'b11111111100000000000001111111111,
            32'b11111111000000000000000111111111,
            32'b11111111000000000000000111111111,
            32'b11111110000000000000000011111111,
            32'b11111110000000000000000011111111,
            32'b11111110000000000000000011111111,
            32'b11111110000000000000000011111111,
            32'b11111110000000000000000011111111,
            32'b11111110000000000000000011111111,
            32'b11111110000000000000000011111111,
            32'b11111110000000000000000011111111,
            32'b11111111000000000000000111111111,
            32'b11111111000000000000000111111111,
            32'b11111111100000000000001111111111,
            32'b11111111110000000000011111111111,
            32'b11111111111000000000111111111111,
            32'b01111111111111111111111111111110,
            32'b00111111111111111111111111111100,
            32'b00011111111111111111111111111000,
            32'b00001111111111111111111111110000,
            32'b00000011111111111111111111000000,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        },

       	{
				32'b00000000000000000000000000000000,
      		32'b00000000000000000000000000000000,
            32'b00000000001111111111000000000000,
            32'b00000000111111111111000000000000,
            32'b00000011111111111111000000000000,
            32'b00001111111111111111000000000000,
            32'b00111111111111111111000000000000,
            32'b11111111111111111111000000000000,
            32'b11111111111111111111000000000000,
            32'b11111111000011111111000000000000,
            32'b11111100000011111111000000000000,
            32'b11111000000011111111000000000000,
            32'b11100000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b00000000000011111111000000000000,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        },

        {
				32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000,
            32'b00000111111111111111111111100000,
            32'b00011111111111111111111111111000,
            32'b00111111111111111111111111111100,
            32'b01111111111111111111111111111110,
            32'b11111111111111111111111111111111,
            32'b11111111100000000000011111111111,
            32'b11111110000000000000001111111111,
            32'b00000000000000000000001111111111,
            32'b00000000000000000000001111111111,
            32'b00000000000000000000011111111110,
            32'b00000000000000000001111111111100,
            32'b00000000000000000111111111111000,
            32'b00000000000000011111111111100000,
            32'b00000000000001111111111110000000,
            32'b00000000000111111111111000000000,
            32'b00000000011111111111100000000000,
            32'b00000001111111111110000000000000,
            32'b00000111111111111000000000000000,
            32'b00011111111111100000000000000000,
            32'b01111111111110000000000000000000,
            32'b11111111111000000000000000000000,
            32'b11111111110000000000000000000000,
            32'b11111111100000000000000000000000,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        },

        {
				32'b00000000000000000000000000000000,
				32'b00000000000000000000000000000000,
            32'b00000011111111111111111000000000,
            32'b00001111111111111111111110000000,
            32'b00111111111111111111111111100000,
            32'b01111111111111111111111111110000,
            32'b11111111111111111111111111111000,
            32'b11111111000000000001111111111100,
            32'b11111100000000000000111111111110,
            32'b00000000000000000000011111111110,
            32'b00000000000000000000011111111110,
            32'b00000000000000000000011111111110,
            32'b00000000000000000000111111111100,
            32'b00000000001111111111111111111000,
            32'b00000000001111111111111111100000,
            32'b00000000001111111111111111100000,
            32'b00000000001111111111111111110000,
            32'b00000000000000000000111111111100,
            32'b00000000000000000000011111111110,
            32'b00000000000000000000001111111110,
            32'b00000000000000000000001111111110,
            32'b00000000000000000000001111111110,
            32'b11111100000000000000011111111100,
            32'b11111111000000000001111111111000,
            32'b11111111111111111111111111110000,
            32'b01111111111111111111111111000000,
            32'b00111111111111111111111100000000,
            32'b00001111111111111111110000000000,
            32'b00000011111111111111000000000000,
            32'b00000000111111111100000000000000,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000,
        },

        {
				32'b00000000000000000000000000000000,
				32'b00000000000000000000000000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000001111111111000000000,
            32'b00000000000111111111111000000000,
            32'b00000000011111111111111000000000,
            32'b00000001111111111111111000000000,
            32'b00000111111111011111111000000000,
            32'b00011111111100011111111000000000,
            32'b01111111110000011111111000000000,
            32'b11111111100000011111111000000000,
            32'b11111111000000011111111000000000,
            32'b11111110000000011111111000000000,
            32'b11111100000000011111111000000000,
            32'b11111000000000011111111000000000,
            32'b11110000000000011111111000000000,
            32'b11100000000000011111111000000000,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b00000000000000011111111000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000000011111111000000000,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        },

        {
				32'b00000000000000000000000000000000,
				32'b00000000000000000000000000000000,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111000000000000000000000000,
            32'b11111111000000000000000000000000,
            32'b11111111000000000000000000000000,
            32'b11111111000000000000000000000000,
            32'b11111111000000000000000000000000,
            32'b11111111000000000000000000000000,
            32'b11111111111111111111111000000000,
            32'b11111111111111111111111110000000,
            32'b11111111111111111111111111100000,
            32'b11111111111111111111111111110000,
            32'b00000000000000000001111111111000,
            32'b00000000000000000000111111111100,
            32'b00000000000000000000011111111110,
            32'b00000000000000000000011111111110,
            32'b00000000000000000000001111111110,
            32'b00000000000000000000001111111110,
            32'b00000000000000000000001111111110,
            32'b00000000000000000000011111111100,
            32'b11111111111111111111111111111000,
            32'b11111111111111111111111111100000,
            32'b11111111111111111111111111000000,
            32'b11111111111111111111111100000000,
            32'b11111111111111111111110000000000,
            32'b00000011111111111111000000000000,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        },

        {
				32'b00000000000000000000000000000000,
				32'b00000000000000000000000000000000,
            32'b00000000111111111111111100000000,
            32'b00000111111111111111111111100000,
            32'b00011111111111111111111111110000,
            32'b00111111111111111111111111111000,
            32'b01111111111000000001111111111100,
            32'b11111111100000000000111111111110,
            32'b11111111000000000000011111111111,
            32'b11111110000000000000001111111111,
            32'b11111110000000000000000111111111,
            32'b11111100000000000000000000000000,
            32'b11111100000000000000000000000000,
            32'b11111100011111111111111000000000,
            32'b11111100111111111111111110000000,
            32'b11111111111111111111111111000000,
            32'b11111111111111111111111111100000,
            32'b11111111111000000011111111110000,
            32'b11111111100000000001111111111000,
            32'b11111111000000000000111111111100,
            32'b11111110000000000000011111111100,
            32'b11111110000000000000011111111100,
            32'b11111110000000000000011111111100,
            32'b11111110000000000000111111111000,
            32'b11111111000000000001111111110000,
            32'b01111111100000000111111111100000,
            32'b00111111111111111111111111000000,
            32'b00011111111111111111111110000000,
            32'b00000111111111111111111000000000,
            32'b00000001111111111111100000000000,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        },

        {
			32'b00000000000000000000000000000000,
			32'b00000000000000000000000000000000,
			32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b11111111111111111111111111111111,
            32'b00000000000000000001111111111110,
            32'b00000000000000000011111111111100,
            32'b00000000000000000111111111111000,
            32'b00000000000000001111111111110000,
            32'b00000000000000011111111111100000,
            32'b00000000000000111111111111000000,
            32'b00000000000001111111111110000000,
            32'b00000000000011111111111100000000,
            32'b00000000000111111111111000000000,
            32'b00000000001111111111110000000000,
            32'b00000000011111111111100000000000,
            32'b00000000111111111111000000000000,
            32'b00000001111111111110000000000000,
            32'b00000011111111111100000000000000,
            32'b00000111111111111000000000000000,
            32'b00001111111111110000000000000000,
            32'b00011111111111100000000000000000,
            32'b00111111111111000000000000000000,
            32'b01111111111110000000000000000000,
            32'b11111111111100000000000000000000,
            32'b11111111111000000000000000000000,
            32'b11111111110000000000000000000000,
            32'b11111111100000000000000000000000,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        },

        {
			32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000,
            32'b00000011111111111111111100000000,
            32'b00001111111111111111111111000000,
            32'b00111111111111111111111111110000,
            32'b01111111111111111111111111111000,
            32'b11111111111000000011111111111100,
            32'b11111111100000000001111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111100000000001111111111100,
            32'b01111111110000000011111111111000,
            32'b00111111111111111111111111110000,
            32'b00011111111111111111111111100000,
            32'b00011111111111111111111111100000,
            32'b00111111111111111111111111110000,
            32'b01111111110000000011111111111000,
            32'b11111111100000000001111111111100,
            32'b11111111000000000000111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111100000000001111111111100,
            32'b11111111110000000011111111111000,
            32'b01111111111111111111111111110000,
            32'b00111111111111111111111111100000,
            32'b00011111111111111111111111000000,
            32'b00000111111111111111111100000000,
            32'b00000001111111111111110000000000,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        },

        {
			32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000,
            32'b00000011111111111111111100000000,
            32'b00001111111111111111111111000000,
            32'b00111111111111111111111111110000,
            32'b01111111111111111111111111111000,
            32'b11111111111000000011111111111100,
            32'b11111111100000000001111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111000000000000111111111110,
            32'b11111111100000000001111111111110,
            32'b11111111110000000111111111111110,
            32'b01111111111111111111111111111110,
            32'b00111111111111111111111111111110,
            32'b00011111111111111111111111111110,
            32'b00001111111111111000111111111110,
            32'b00000000000000000000111111111110,
            32'b00000000000000000000111111111110,
            32'b00000000000000000000111111111110,
            32'b00000000000000000000111111111100,
            32'b11111100000000000001111111111000,
            32'b11111111000000000111111111110000,
            32'b11111111111111111111111111100000,
            32'b01111111111111111111111111000000,
            32'b00111111111111111111111100000000,
            32'b00001111111111111111110000000000,
            32'b00000011111111111111000000000000,
            32'b00000000111111111100000000000000,
            32'b00000000000000000000000000000000,
            32'b00000000000000000000000000000000
        }
};


 

logic [0:1] [0:31] [0:31] levelLabel  = {
	{
		32'b	00000000000000000000000000000000,
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111110000000000000000000000, 
		32'b	11111111111111111111111111111111,
		32'b	11111111111111111111111111111111,
		32'b	11111111111111111111111111111111,
		32'b	11111111111111111111111111111111,
		32'b	11111111111111111111111111111111,
		32'b	11111111111111111111111111111111,
		32'b	11111111111111111111111111111111,
	},
	{
		32'b    00000000000000000000000000000000,
		32'b    00000000000000000000000000000000,
		32'b    00000000000000000000000000000000,
		32'b    00000000000000000000000000000000,
		32'b    00000000000000000000000000000000,
		32'b    00000000000000000000000000000000,
		32'b    00000000000000000000000000000000,
		32'b	00000000000000000000000000000000,
		32'b 	00000000000000000000000000000000,
		32'b 	00000000000000000000000000000000,
		32'b 	00000000000000000000000000000000,
		32'b 	00000000000000000000000000000000,
		32'b 	00000000000000000000000000000000,
		32'b    11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b	11111000000000000011111000000000,
		32'b 	11111000000000000011111000000000,
		32'b 	01111100000000000111110000000000,
		32'b    00111110000000001111100111111100,
		32'b	00011111000000011111001111111110,
		32'b	00001111100000111110011111111111,
		32'b	00000111110001111100011111111111,
		32'b	00000011111011111000001111111110,
		32'b	00000011111111110000000111111100,
	}
};
 
logic [0:31] [0:31] [7:0]  object_colors  = {
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'he4,8'he4,8'he4,8'hFF,8'hFF,8'he4,8'he4,8'he4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h20,8'hed,8'hed,8'he4,8'he4,8'h20,8'h20,8'he4,8'he4,8'he4,8'he4,8'h20,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'hed,8'hFE,8'hFE,8'hed,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'hed,8'hFE,8'hFE,8'hed,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'he4,8'hed,8'hed,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'he0,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'ha0,8'hc0,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hc0,8'ha0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'he0,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'ha0,8'hc0,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hc0,8'ha0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'he0,8'he4,8'he4,8'he0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'ha0,8'hc0,8'he4,8'he4,8'hc0,8'ha0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'ha0,8'ha0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
	{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF}
};

// assign _LSB  = offsetY[4:0] ; // get lower 5 bits 
// assign offsetY_MSB  = offsetY[8:5] ; // get higher 4 bits 
// assign offsetX_LSB  = offsetX[4:0] ; 
// assign offsetX_MSB  = offsetX[8:5] ; 

// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask  <=  MazeDefaultBitMapMask ;  //  copy default tabel 
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
		drawingRequest <= 1'b0;
		
		if (InsideRectangle == 1'b1 )	
			begin 
				// RGBout <= text_color;
		   	case (MazeBitMapMask[offsetX[8:5]])
					 4'h0 : RGBout <= TRANSPARENT_ENCODING ;
					 4'hA : begin 
							drawingRequest <= levelLabel[0][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'hB : begin 
							drawingRequest <= levelLabel[1][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h8 : begin 
							drawingRequest <= number_bitmap[level+1][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h9 : begin 
							drawingRequest <= number_bitmap[birdsLeft][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'hC : begin 
							drawingRequest <= (object_colors[offsetY[4:0]][offsetX[4:0]] != TRANSPARENT_ENCODING) ? 1'b1 : 1'b0;
							RGBout <= object_colors[offsetY[4:0]][offsetX[4:0]];
					 end
					 4'h3 : begin 
							drawingRequest <= number_bitmap[0][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h4 : begin 
							drawingRequest <= number_bitmap[score[3:0]][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h5 : begin 
							drawingRequest <= number_bitmap[score[7:4]][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h6 : begin 
							drawingRequest <= number_bitmap[score[11:8]][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					//  4'h2 : RGBout <= object_colors[2'h1][offsetY[4:0]][offsetX[4:0]] ; 
					 default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
			end 
 
	end 
end
//
////==----------------------------------------------------------------------------------------------------------------=
//// decide if to draw the pixel or not 
//assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

