// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	StatsDisplayBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,// offset from top left  position 
					input logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic [3:0] level,
					input logic [3:0] birdsLeft,
					input logic [11:0] score,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 

parameter  logic	[7:0] text_color = 8'h00 ; //set the color of the digit 


logic [0:15] [3:0]  MazeBitMapMask ;  

// A - level number (based on input)
// C - number of birds left (based on input)
// 1 - level label
// 2 - heart label
// 3 - score digit (based on input)
// 4 - score digit (based on input)
// 5 - score digit (based on input)
// 6 - score digit (based on input)
logic [0:15] [3:0]  MazeDefaultBitMapMask= 64'h01A000C200065430;
 
 
bit [0:9] [0:31] [0:31] number_bitmap  = {

{32'b	00000000000000000000000000000000,
32'b	00000000001111111100000000000000,
32'b	00000011111111111111110000000000,
32'b	00001111111111111111111100000000,
32'b	00011111111111111111111110000000,
32'b	00111111100000000001111111000000,
32'b	01111111000000000000011111100000,
32'b	01111110000000000000001111110000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	01111110000000000000001111110000,
32'b	01111111000000000000011111100000,
32'b	00111111100000000001111111000000,
32'b	00011111111111111111111110000000,
32'b	00001111111111111111111100000000,
32'b	00000011111111111111110000000000,
32'b	00000000001111111100000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000
},
																	
{32'b	00000000000001111110000000000000,
32'b	00000000000011111110000000000000,
32'b	00000000000111111110000000000000,
32'b	00000000001111111110000000000000,
32'b	00000000011111111110000000000000,
32'b	00000000111111111110000000000000,
32'b	00000001111111011110000000000000,
32'b	00000011111100011110000000000000,
32'b	00000111110000011110000000000000,
32'b	00001111100000011110000000000000,
32'b	00011111000000011110000000000000,
32'b	00111110000000011110000000000000,
32'b	01111100000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	00000000000000011110000000000000,
32'b	01111111111111111111111111111110,
32'b	01111111111111111111111111111110,
32'b	01111111111111111111111111111110,
32'b	01111111111111111111111111111110,
32'b	01111111111111111111111111111110,
},

																	

{
32'b	00000000000000000000000000000000,
32'b	00000000001111111100000000000000,
32'b	00000011111111111111110000000000,
32'b	00001111111111111111111100000000,
32'b	00011111111111111111111110000000,
32'b	00111111100000000001111111000000,
32'b	01111111000000000000011111100000,
32'b	01111110000000000000001111110000,
32'b	11111100000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	00000000000000000000000111111000,
32'b	00000000000000000000001111110000,
32'b	00000000000000000000011111100000,
32'b	00000000000000000000111111000000,
32'b	00000000000000000001111110000000,
32'b	00000000000000000011111100000000,
32'b	00000000000000001111111000000000,
32'b	00000000000000011111110000000000,
32'b	00000000000000111111100000000000,
32'b	00000000000001111111000000000000,
32'b	00000000000011111110000000000000,
32'b	00000000000111111100000000000000,
32'b	00000000001111111000000000000000,
32'b	00000000011111110000000000000000,
32'b	00000000111111100000000000000000,
32'b	00000001111111000000000000000000,
32'b	00000011111110000000000000000000,
32'b	00000111111111111111111111111110,
32'b	00001111111111111111111111111110,
32'b	00011111111111111111111111111110,
32'b	00111111111111111111111111111110,
32'b	01111111111111111111111111111110,
},

																	
{32'b	00000000001111111100000000000000,
32'b	00000011111111111111110000000000,
32'b	00001111111111111111111100000000,
32'b	00011111111111111111111110000000,
32'b	00111111100000000001111111000000,
32'b	01111111000000000000011111100000,
32'b	01111110000000000000001111110000,
32'b	11111100000000000000000111111000,
32'b	00000000000000000000000111111000,
32'b	00000000000000000000001111110000,
32'b	00000000000000000000111111100000,
32'b	00000000000011111111111111000000,
32'b	00000000000011111111111100000000,
32'b	00000000000011111111111111000000,
32'b	00000000000000000000111111100000,
32'b	00000000000000000000001111110000,
32'b	00000000000000000000000111111000,
32'b	00000000000000000000000111111000,
32'b	11111100000000000000000111111000,
32'b	01111110000000000000001111110000,
32'b	01111111000000000000011111100000,
32'b	00111111100000000001111111000000,
32'b	00011111111111111111111110000000,
32'b	00001111111111111111111100000000,
32'b	00000011111111111111110000000000,
32'b	00000000001111111100000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000},

																	
{32'b	00000000000000000001111000000000,
32'b	00000000000000000001111000000000,
32'b	00000000000000000011111000000000,
32'b	00000000000000000111111000000000,
32'b	00000000000000001111111000000000,
32'b	00000000000000011111111000000000,
32'b	00000000000000111111111000000000,
32'b	00000000000001111111111000000000,
32'b	00000000000011111011111000000000,
32'b	00000000000111110011111000000000,
32'b	00000000001111100011111000000000,
32'b	00000000011111000011111000000000,
32'b	00000000111110000011111000000000,
32'b	00000001111100000011111000000000,
32'b	00000011111000000011111000000000,
32'b	00000111110000000011111000000000,
32'b	00001111111111111111111111111110,
32'b	00001111111111111111111111111110,
32'b	00001111111111111111111111111110,
32'b	00001111111111111111111111111110,
32'b	00000000000000000011111000000000,
32'b	00000000000000000011111000000000,
32'b	00000000000000000011111000000000,
32'b	00000000000000000011111000000000,
32'b	00000000000000000011111000000000,
32'b	00000000000000000011111000000000,
32'b	00000000000000000011111000000000,
32'b	00000000000000000011111000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000},

																	
{32'b	00000011111111111111111111111100,
32'b	00000011111111111111111111111100,
32'b	00000011111111111111111111111100,
32'b	00000011111111111111111111111100,
32'b	00000011111110000000000000000000,
32'b	00000011111110000000000000000000,
32'b	00000011111110000000000000000000,
32'b	00000011111110000000000000000000,
32'b	00000011111111111111111111000000,
32'b	00000011111111111111111111110000,
32'b	00000011111111111111111111111000,
32'b	00000011111111111111111111111100,
32'b	00000000000000000000011111111100,
32'b	00000000000000000000000111111100,
32'b	00000000000000000000000011111100,
32'b	00000000000000000000000011111100,
32'b	11111100000000000000000011111100,
32'b	11111100000000000000000011111100,
32'b	11111100000000000000000011111100,
32'b	11111110000000000000000111111100,
32'b	01111111000000000000011111111100,
32'b	01111111110000000011111111111000,
32'b	00111111111111111111111111111000,
32'b	00011111111111111111111111110000,
32'b	00001111111111111111111111100000,
32'b	00000011111111111111111110000000,
32'b	00000000001111111111111000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000},

																	
{32'b	00000000000000000011111111000000,
32'b	00000000001111111111111111110000,
32'b	00000000111111111111111111111000,
32'b	00000001111111111111111111111100,
32'b	00000011111111111111110000000000,
32'b	00000111111111000000000000000000,
32'b	00001111111100000000000000000000,
32'b	00011111110000000000000000000000,
32'b	00111111100000000000000000000000,
32'b	01111111000000000000000000000000,
32'b	11111111111111111111111111000000,
32'b	11111111111111111111111111110000,
32'b	11111111111111111111111111111000,
32'b	11111111111111111111111111111100,
32'b	11111111000000000000111111111100,
32'b	11111110000000000000001111111100,
32'b	11111100000000000000000111111100,
32'b	11111100000000000000000111111100,
32'b	11111100000000000000000111111100,
32'b	01111110000000000000001111111100,
32'b	01111111000000000000111111111000,
32'b	00111111110000000011111111111000,
32'b	00011111111111111111111111110000,
32'b	00001111111111111111111111100000,
32'b	00000111111111111111111110000000,
32'b	00000000111111111111111100000000,
32'b	00000000000111111111110000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000},

																	
{32'b	01111111111111111111111111111110,
32'b	01111111111111111111111111111110,
32'b	01111111111111111111111111111110,
32'b	01111111111111111111111111111110,
32'b	00000000000000000001111111000000,
32'b	00000000000000000011111110000000,
32'b	00000000000000000011111100000000,
32'b	00000000000000000111111100000000,
32'b	00000000000000001111111000000000,
32'b	00000000000000011111110000000000,
32'b	00000000000000111111100000000000,
32'b	00000000000001111111000000000000,
32'b	00000000000011111110000000000000,
32'b	00000000000111111100000000000000,
32'b	00000000001111111000000000000000,
32'b	00000000011111110000000000000000,
32'b	00000000111111100000000000000000,
32'b	00000001111111000000000000000000,
32'b	00000011111110000000000000000000,
32'b	00000111111100000000000000000000,
32'b	00001111111000000000000000000000,
32'b	00011111110000000000000000000000,
32'b	00111111100000000000000000000000,
32'b	01111111000000000000000000000000,
32'b	11111110000000000000000000000000,
32'b	11111100000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000},

																	
{32'b	00000000001111111111100000000000,
32'b	00000001111111111111111000000000,
32'b	00000111111111111111111110000000,
32'b	00001111111111111111111111000000,
32'b	00011111110000000000111111100000,
32'b	00111111100000000000011111110000,
32'b	01111111000000000000001111111000,
32'b	01111110000000000000000111111000,
32'b	01111110000000000000000111111000,
32'b	01111110000000000000000111111000,
32'b	00111111000000000000001111110000,
32'b	00111111100000000000011111100000,
32'b	00011111111000000001111111000000,
32'b	00001111111110000111111110000000,
32'b	00000111111111111111111100000000,
32'b	00000011111111111111111000000000,
32'b	00000111111111111111111100000000,
32'b	00011111111000000001111111100000,
32'b	00111111100000000000011111110000,
32'b	01111111000000000000001111111000,
32'b	11111110000000000000000111111100,
32'b	11111110000000000000000111111100,
32'b	11111110000000000000000111111100,
32'b	01111111000000000000001111111000,
32'b	01111111100000000000011111111000,
32'b	00111111111100000001111111110000,
32'b	00011111111111111111111111100000,
32'b	00001111111111111111111111000000,
32'b	00000011111111111111111100000000,
32'b	00000000111111111111110000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000},
															
{32'b	00000000001111111111100000000000,
32'b	00000001111111111111111000000000,
32'b	00000111111111111111111110000000,
32'b	00001111111111111111111111000000,
32'b	00011111111000000000111111100000,
32'b	00111111100000000000011111110000,
32'b	01111111000000000000001111111000,
32'b	01111110000000000000000111111000,
32'b	11111110000000000000000111111100,
32'b	11111110000000000000000111111100,
32'b	11111110000000000000000111111100,
32'b	11111110000000000000000111111100,
32'b	01111111000000000000001111111100,
32'b	00111111100000000000011111111100,
32'b	00011111111111111111111111111000,
32'b	00001111111111111111111111111000,
32'b	00000111111111111111111111110000,
32'b	00000001111111111111111111000000,
32'b	00000000000000000000011111100000,
32'b	00000000000000000000001111110000,
32'b	00000000000000000000000111110000,
32'b	00000000000000000000001111100000,
32'b	00000000000000000000011111100000,
32'b	00000000000000000011111111000000,
32'b	00000011111111111111111110000000,
32'b	00000111111111111111111100000000,
32'b	00001111111111111111111000000000,
32'b	00001111111111111111110000000000,
32'b	00000011111111111110000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000,
32'b	00000000000000000000000000000000},
} ; 


 

logic [0:31] [0:31] levelLabel  = {
	32'b	11111000000000000000000000000000, 
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000000000000000000000000000,
	32'b	11111000111100000000000000011110,
	32'b	11111000011110000000000000111100,
	32'b	11111000001111000000000001111000,
	32'b	11111000000111100000000011110000,
	32'b	11111000000011110000000111100000,
	32'b	11111000000001111000001111011100,
	32'b	11111111111100111100011110110110,
	32'b	11111111111100011110111101100011,
	32'b	11111111111100001111111000110110,
	32'b	11111111111100000111110000011100,
};
 
logic [0:31] [0:31] [7:0]  object_colors  = {
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'hAC, 8'hCD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'hC1, 8'hC1, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB0, 8'h78, 8'h3C, 8'h1C, 8'h55, 8'hCD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA9, 8'h62, 8'h87, 8'hC7, 8'hE7, 8'hE3, 8'hC2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'h9C, 8'h7C, 8'h3C, 8'h3C, 8'h1D, 8'h39, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hA9, 8'h26, 8'h47, 8'h87, 8'hC3, 8'hE7, 8'hE7, 8'hE7, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD4, 8'hBC, 8'h7C, 8'h3C, 8'h1C, 8'h3D, 8'h1E, 8'h3A, 8'hAD, 8'hFF, 8'hCE, 8'h26, 8'h27, 8'h67, 8'h83, 8'hC7, 8'hE7, 8'hE7, 8'hE3, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD8, 8'hBC, 8'h7C, 8'h5C, 8'h3C, 8'h1D, 8'h3E, 8'h1E, 8'h3A, 8'hCD, 8'h4E, 8'h0B, 8'h27, 8'h47, 8'h87, 8'hA3, 8'hE7, 8'hE7, 8'hE7, 8'hE6, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hDC, 8'hBC, 8'h7C, 8'h5C, 8'h3C, 8'h3D, 8'h1D, 8'h1E, 8'h1F, 8'h52, 8'h2F, 8'h0B, 8'h27, 8'h47, 8'h87, 8'hA7, 8'hE7, 8'hE7, 8'hE7, 8'hE7, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hFC, 8'hBC, 8'h9C, 8'h5C, 8'h3C, 8'h1D, 8'h3D, 8'h1E, 8'h1F, 8'h1B, 8'h13, 8'h0B, 8'h27, 8'h47, 8'h86, 8'hA6, 8'hE7, 8'hE7, 8'hE7, 8'hE3, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hFC, 8'hBC, 8'h9C, 8'h5C, 8'h3C, 8'h3D, 8'h1D, 8'h1E, 8'h1F, 8'h1B, 8'h13, 8'h0F, 8'h27, 8'h47, 8'hA0, 8'hA0, 8'hC6, 8'hE7, 8'hE7, 8'hE7, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hFC, 8'hBC, 8'h9C, 8'h5C, 8'h3C, 8'h1D, 8'h3D, 8'h3A, 8'h3E, 8'h3B, 8'h13, 8'h0F, 8'h07, 8'h47, 8'hA0, 8'hC0, 8'hC6, 8'hE7, 8'hE7, 8'hE3, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hFC, 8'hDC, 8'h9C, 8'h5C, 8'h3C, 8'h1C, 8'h68, 8'h6D, 8'h56, 8'h85, 8'h4E, 8'h0F, 8'h07, 8'h27, 8'h81, 8'hA1, 8'hC7, 8'hE7, 8'hE7, 8'hE7, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hFC, 8'hDC, 8'h9C, 8'h7C, 8'h3C, 8'h6C, 8'hC0, 8'h84, 8'h51, 8'hC0, 8'h85, 8'h0F, 8'h0B, 8'h27, 8'h66, 8'h86, 8'hA1, 8'hC2, 8'hE7, 8'hE7, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hF8, 8'hDC, 8'h9C, 8'h7C, 8'h3C, 8'h50, 8'hC0, 8'hA4, 8'h56, 8'hC0, 8'h69, 8'h2E, 8'h26, 8'h46, 8'h81, 8'h82, 8'hA0, 8'hC1, 8'hE7, 8'hE3, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hF8, 8'hDC, 8'hBC, 8'h7C, 8'h74, 8'h54, 8'h84, 8'h89, 8'h3E, 8'h6D, 8'h4E, 8'hA0, 8'h65, 8'h61, 8'hA0, 8'hA0, 8'hC0, 8'hC1, 8'hC7, 8'hE7, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hDC, 8'hBC, 8'h94, 8'hA0, 8'hA0, 8'h51, 8'h39, 8'h1E, 8'h1F, 8'h69, 8'hC0, 8'h81, 8'h80, 8'hC0, 8'hC0, 8'hC0, 8'hC1, 8'hC7, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hFC, 8'hBC, 8'h98, 8'hA0, 8'hA0, 8'h88, 8'h1D, 8'h3A, 8'h4D, 8'h69, 8'hC0, 8'h85, 8'h80, 8'hC0, 8'hC0, 8'hC0, 8'hC1, 8'hC6, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hFC, 8'hAC, 8'h88, 8'hC0, 8'hC0, 8'h84, 8'h3D, 8'h55, 8'hC0, 8'h69, 8'h89, 8'h66, 8'h80, 8'hC0, 8'hC0, 8'hC0, 8'hC1, 8'hC3, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hD8, 8'hA0, 8'hC0, 8'hC0, 8'hC0, 8'h84, 8'h51, 8'h69, 8'hC0, 8'h69, 8'h17, 8'h2F, 8'h65, 8'hA0, 8'hC0, 8'hC0, 8'hA1, 8'hC2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD0, 8'hC4, 8'hC0, 8'hC0, 8'hC0, 8'h84, 8'h84, 8'hC0, 8'hC0, 8'h89, 8'h17, 8'h0F, 8'h26, 8'h80, 8'hC0, 8'hC0, 8'hC6, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hC8, 8'hC0, 8'hC0, 8'hC0, 8'h88, 8'h88, 8'hC0, 8'hC0, 8'h89, 8'h33, 8'h2E, 8'h45, 8'h61, 8'hA0, 8'hC0, 8'hC2, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAC, 8'hC4, 8'hC0, 8'hC0, 8'h8C, 8'h70, 8'hC0, 8'hC0, 8'h89, 8'h69, 8'h65, 8'hA0, 8'h81, 8'h66, 8'hA1, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'h90, 8'hC0, 8'hC0, 8'h6C, 8'h1D, 8'h6D, 8'hA4, 8'h6D, 8'hA4, 8'hC0, 8'hC0, 8'h80, 8'h47, 8'h83, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h94, 8'h74, 8'h88, 8'h54, 8'h1D, 8'h1E, 8'h3E, 8'h3A, 8'h85, 8'hC0, 8'hC0, 8'h81, 8'h47, 8'h82, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'h7C, 8'h5C, 8'h1C, 8'h1D, 8'h3D, 8'h69, 8'h6D, 8'h4E, 8'hA0, 8'hC0, 8'h61, 8'h43, 8'hAA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h94, 8'h5C, 8'h3C, 8'h1D, 8'h39, 8'hC0, 8'h89, 8'h37, 8'h84, 8'hC0, 8'h46, 8'h66, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'h58, 8'h3C, 8'h1D, 8'h3D, 8'hA4, 8'h6D, 8'h1B, 8'h52, 8'h85, 8'h27, 8'hAA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h90, 8'h3C, 8'h1D, 8'h1D, 8'h3A, 8'h3A, 8'h1B, 8'h13, 8'h0F, 8'h66, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h54, 8'h1C, 8'h3D, 8'h1E, 8'h1E, 8'h3B, 8'h17, 8'h2A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB1, 8'h3C, 8'h1D, 8'h1E, 8'h1E, 8'h1B, 8'h17, 8'h8D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h70, 8'h1D, 8'h3E, 8'h3E, 8'h1F, 8'h6E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h1E, 8'h1E, 8'h56, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'h39, 8'h3A, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
	{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF }
};

// assign _LSB  = offsetY[4:0] ; // get lower 5 bits 
// assign offsetY_MSB  = offsetY[8:5] ; // get higher 4 bits 
// assign offsetX_LSB  = offsetX[4:0] ; 
// assign offsetX_MSB  = offsetX[8:5] ; 

// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask  <=  MazeDefaultBitMapMask ;  //  copy default tabel 
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
		drawingRequest <= 1'b0;
		
		if (InsideRectangle == 1'b1 )	
			begin 
				// RGBout <= text_color;
		   	case (MazeBitMapMask[offsetX[8:5]])
					 4'h0 : RGBout <= TRANSPARENT_ENCODING ;
					 4'h1 : begin 
							drawingRequest <= levelLabel[offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'hA : begin 
							drawingRequest <= number_bitmap[level+1][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'hC : begin 
							drawingRequest <= number_bitmap[birdsLeft][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h2 : begin 
							drawingRequest <= (object_colors[offsetY[4:0]][offsetX[4:0]] != TRANSPARENT_ENCODING) ? 1'b1 : 1'b0;
							RGBout <= object_colors[offsetY[4:0]][offsetX[4:0]];
					 end
					 4'h3 : begin 
							drawingRequest <= number_bitmap[0][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h4 : begin 
							drawingRequest <= number_bitmap[score[3:0]][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h5 : begin 
							drawingRequest <= number_bitmap[score[7:4]][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					 4'h5 : begin 
							drawingRequest <= number_bitmap[score[11:8]][offsetY[4:0]][offsetX[4:0]];
							RGBout <= text_color;
					 end
					//  4'h2 : RGBout <= object_colors[2'h1][offsetY[4:0]][offsetX[4:0]] ; 
					 default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
			end 
 
	end 
end
//
////==----------------------------------------------------------------------------------------------------------------=
//// decide if to draw the pixel or not 
//assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

