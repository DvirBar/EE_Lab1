// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  2023  
// (c) Technion IIT, Department of Electrical Engineering 2023 



module	StatsDisplayBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic random_hart,
					
//------------------------input collision smiley and hart -student to complete functionality					
					input smiley_hart_collision,
			

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 


logic [0:15] [0:15] [3:0]  MazeBitMapMask ;  

logic [0:15] [0:15] [3:0]  MazeDefaultBitMapMask= // defult table to load on reset 
{{64'h0001110000011100},
 {64'h0010002102100010},
 {64'h0010000010000010},
 {64'h0001000000000100},
 {64'h0001000000000100},
 {64'h0000100000001000},
 {64'h0000010000010000},
 {64'h0000001000100000},
 {64'h0000000101000000},
 {64'h0000000010000000},
 {64'h0000000000000000},
 {64'h0002000000002000},
 {64'h0000000000000000},
 {64'h0000000000000000},
 {64'h0000000000000000},
 {64'h0000000000000000}};
 
 
bit [0:15] [0:31] [0:15] number_bitmap  = {

{16'b	0000001111100000,
16'b	0000111111111000,
16'b	0000111111111000,
16'b	0001111111111100,
16'b	0011111001111100,
16'b	0011100000111110,
16'b	0111100000011110,
16'b	0111100000011110,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000011110,
16'b	1111100000011110,
16'b	0111110000111110,
16'b	0111110000111100,
16'b	0011111001111100,
16'b	0011111111111000,
16'b	0001111111111000,
16'b	0000111111110000,
16'b	0000011111000000},


																	
{16'b	0000000011100000,
16'b	0000000111100000,
16'b	0000011111100000,
16'b	0000111111100000,
16'b	0001111111100000,
16'b	0011111111100000,
16'b	0111111011100000,
16'b	0111100011100000,
16'b	0111000011100000,
16'b	0010000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111111},
																	
{16'b	0000111111100000,
16'b	0001111111110000,
16'b	0111111111111000,
16'b	1111111111111000,
16'b	1111110011111100,
16'b	1111000011111100,
16'b	1110000001111110,
16'b	0000000000111110,
16'b	0000000000111110,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000001111100,
16'b	0000000001111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011110000,
16'b	0000000011100000,
16'b	0000000111000000,
16'b	0000001111000000,
16'b	0000011110000000,
16'b	0000111100000000,
16'b	0001111100000000,
16'b	0001111100000000,
16'b	0011111000000000,
16'b	0111110000000001,
16'b	1111100000000011,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111},
																	
{16'b	0000111111100000,
16'b	0001111111111000,
16'b	0111111111111000,
16'b	1111111111111000,
16'b	1111110011111100,
16'b	1111000001111100,
16'b	1110000001111100,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000000111100,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0001111111110000,
16'b	0001111111000000,
16'b	0001111111111000,
16'b	0001111111111000,
16'b	0000000011111100,
16'b	0000000001111110,
16'b	0000000000111111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000111111,
16'b	1110000001111110,
16'b	1111100011111110,
16'b	1111111111111100,
16'b	1111111111111000,
16'b	0111111111111000,
16'b	0001111111000000},
																	
{16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000111111000,
16'b	0000001111111000,
16'b	0000001101111000,
16'b	0000011101111000,
16'b	0000011101111000,
16'b	0000111101111000,
16'b	0001111101111000,
16'b	0001111101111000,
16'b	0001111001111000,
16'b	0011111001111000,
16'b	0011110001111000,
16'b	0111100001111000,
16'b	0111100001111000,
16'b	1111000001111000,
16'b	1110000001111000,
16'b	1110000001111000,
16'b	1110000001111000,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000011111100},
																	
{16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111110,
16'b	0111111111111100,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111111111100000,
16'b	0111111111111000,
16'b	0111111111111000,
16'b	0111111111111100,
16'b	0010000011111110,
16'b	0000000001111110,
16'b	0000000000111111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	1000000000111110,
16'b	1100000001111110,
16'b	1111100011111100,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	0001111111000000},
																	
{16'b	0000000111111100,
16'b	0000011111111110,
16'b	0000111111111110,
16'b	0001111111111111,
16'b	0001111100001111,
16'b	0011111100000001,
16'b	0011111000000000,
16'b	0111110000000000,
16'b	0111100000000000,
16'b	1111100000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111001111111000,
16'b	1111111111111100,
16'b	1111111111111110,
16'b	1111111111111111,
16'b	1111111101111111,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111100000001111,
16'b	1111100000001111,
16'b	0111110000011111,
16'b	0111111101111110,
16'b	0011111111111110,
16'b	0001111111111100,
16'b	0001111111111000,
16'b	0000011111100000},
																	
{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1100000000001111,
16'b	1000000000011111,
16'b	0000000000011111,
16'b	0000000000011110,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000001111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011110000,
16'b	0000000011110000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000111100000,
16'b	0000000111100000,
16'b	0000001111000000,
16'b	0000001111000000,
16'b	0000011110000000,
16'b	0000011110000000,
16'b	0000111110000000,
16'b	0000111100000000,
16'b	0000111100000000,
16'b	0001111100000000,
16'b	0001111100000000,
16'b	0001111100000000},
																	
{16'b	0000111111110000,
16'b	0001111111111000,
16'b	0011111111111100,
16'b	0111111111111110,
16'b	0111111011111110,
16'b	1111100000111111,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111100000011110,
16'b	0111110000111110,
16'b	0111111001111100,
16'b	0011111111111000,
16'b	0001111111111000,
16'b	0000111111100000,
16'b	0000111111110000,
16'b	0001111111111000,
16'b	0011111111111100,
16'b	0111111001111110,
16'b	1111100000111111,
16'b	1111000000001111,
16'b	1110000000001111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1111000000001111,
16'b	1111100000011111,
16'b	1111111001111111,
16'b	1111111111111110,
16'b	0111111111111110,
16'b	0011111111111000,
16'b	0001111111110000},
																	
{16'b	0000111111100000,
16'b	0001111111111000,
16'b	0011111111111000,
16'b	0111111111111100,
16'b	1111111011111100,
16'b	1111100000111110,
16'b	1111000000011110,
16'b	1111000000011111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1111000000001111,
16'b	1111100000011111,
16'b	1111111011111111,
16'b	1111111111111111,
16'b	0111111111111111,
16'b	0011111111111111,
16'b	0001111111001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000011110,
16'b	0000000000011110,
16'b	0000000000111110,
16'b	0000000001111100,
16'b	1000000011111100,
16'b	1111000011111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	1111111111100000,
16'b	0011111100000000},

{16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000111111110000,
16'b	0000110000111000,
16'b	0000110000111000,
16'b	0000110000111000,
16'b	0001110000111100,
16'b	0001100000011100,
16'b	0011100000011100,
16'b	0011000000001100,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1111000000001111},


{16'b	1111111111110000,
16'b	1111111111111000,
16'b	1111111111111100,
16'b	1111111111111110,
16'b	0111000011111110,
16'b	0111000000111111,
16'b	0111000000011111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000011110,
16'b	0111000000111110,
16'b	0111000001111100,
16'b	0111111111111000,
16'b	0111111111111000,
16'b	0111111111100000,
16'b	0111111111110000,
16'b	0111111111111000,
16'b	0111111111111100,
16'b	0111000001111110,
16'b	0111000000111111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000000111,
16'b	0111000000000111,
16'b	0111000000001111,
16'b	0111000000011111,
16'b	0111000001111111,
16'b	1111111111111110,
16'b	1111111111111110,
16'b	1111111111111000,
16'b	1111111111110000},

{16'b	0000001111111000,
16'b	0000111111111100,
16'b	0000111111111110,
16'b	0001111111111111,
16'b	0011111001000011,
16'b	0011100000000001,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	1111100000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111100000000000,
16'b	0111110000000000,
16'b	0111110000000001,
16'b	0011111001000011,
16'b	0011111111111111,
16'b	0001111111111110,
16'b	0000111111111100,
16'b	0000011111111000},


{16'b	1111111111100000,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111111100,
16'b	0111000001111100,
16'b	0111000000111110,
16'b	0111000000011110,
16'b	0111000000011110,
16'b	0111000000011111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000011110,
16'b	0111000000011110,
16'b	0111000000111110,
16'b	0111000000111100,
16'b	0111000001111100,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	1111111111000000},

{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000011,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000001,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000001,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000001000011,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111},

{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000011,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000001,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000001,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000}


} ; 


 

 logic [1:0] [0:31] [0:31] [7:0]  object_colors  = {
	 {16'b	0000001111100000,
	16'b	0000111111111000,
	16'b	0000111111111000,
	16'b	0001111111111100,
	16'b	0011111001111100,
	16'b	0011100000111110,
	16'b	0111100000011110,
	16'b	0111100000011110,
	16'b	1111100000011111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000011110,
	16'b	1111100000011110,
	16'b	0111110000111110,
	16'b	0111110000111100,
	16'b	0011111001111100,
	16'b	0011111111111000,
	16'b	0001111111111000,
	16'b	0000111111110000,
	16'b	0000011111000000},


																		
	{16'b	0000000011100000,
	16'b	0000000111100000,
	16'b	0000011111100000,
	16'b	0000111111100000,
	16'b	0001111111100000,
	16'b	0011111111100000,
	16'b	0111111011100000,
	16'b	0111100011100000,
	16'b	0111000011100000,
	16'b	0010000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0111111111111111,
	16'b	0111111111111111,
	16'b	0111111111111111,
	16'b	0111111111111111},
																		
	{16'b	0000111111100000,
	16'b	0001111111110000,
	16'b	0111111111111000,
	16'b	1111111111111000,
	16'b	1111110011111100,
	16'b	1111000011111100,
	16'b	1110000001111110,
	16'b	0000000000111110,
	16'b	0000000000111110,
	16'b	0000000000111110,
	16'b	0000000000111100,
	16'b	0000000001111100,
	16'b	0000000001111100,
	16'b	0000000001111000,
	16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0000000011110000,
	16'b	0000000011100000,
	16'b	0000000111000000,
	16'b	0000001111000000,
	16'b	0000011110000000,
	16'b	0000111100000000,
	16'b	0001111100000000,
	16'b	0001111100000000,
	16'b	0011111000000000,
	16'b	0111110000000001,
	16'b	1111100000000011,
	16'b	1111111111111111,
	16'b	1111111111111111,
	16'b	1111111111111111,
	16'b	1111111111111111},
																		
	{16'b	0000111111100000,
	16'b	0001111111111000,
	16'b	0111111111111000,
	16'b	1111111111111000,
	16'b	1111110011111100,
	16'b	1111000001111100,
	16'b	1110000001111100,
	16'b	0000000000111110,
	16'b	0000000000111100,
	16'b	0000000000111100,
	16'b	0000000000111100,
	16'b	0000000001111100,
	16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0001111111110000,
	16'b	0001111111000000,
	16'b	0001111111111000,
	16'b	0001111111111000,
	16'b	0000000011111100,
	16'b	0000000001111110,
	16'b	0000000000111111,
	16'b	0000000000011111,
	16'b	0000000000011111,
	16'b	0000000000011111,
	16'b	0000000000011111,
	16'b	0000000000111111,
	16'b	1110000001111110,
	16'b	1111100011111110,
	16'b	1111111111111100,
	16'b	1111111111111000,
	16'b	0111111111111000,
	16'b	0001111111000000},
																		
	{16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0000000111111000,
	16'b	0000001111111000,
	16'b	0000001101111000,
	16'b	0000011101111000,
	16'b	0000011101111000,
	16'b	0000111101111000,
	16'b	0001111101111000,
	16'b	0001111101111000,
	16'b	0001111001111000,
	16'b	0011111001111000,
	16'b	0011110001111000,
	16'b	0111100001111000,
	16'b	0111100001111000,
	16'b	1111000001111000,
	16'b	1110000001111000,
	16'b	1110000001111000,
	16'b	1110000001111000,
	16'b	1111111111111111,
	16'b	1111111111111111,
	16'b	1111111111111111,
	16'b	0000000001111000,
	16'b	0000000001111000,
	16'b	0000000001111000,
	16'b	0000000001111000,
	16'b	0000000001111000,
	16'b	0000000001111000,
	16'b	0000000001111000,
	16'b	0000000011111100},
																		
	{16'b	0111111111111111,
	16'b	0111111111111111,
	16'b	0111111111111110,
	16'b	0111111111111100,
	16'b	0111100000000000,
	16'b	0111100000000000,
	16'b	0111100000000000,
	16'b	0111100000000000,
	16'b	0111100000000000,
	16'b	0111100000000000,
	16'b	0111100000000000,
	16'b	0111111111100000,
	16'b	0111111111111000,
	16'b	0111111111111000,
	16'b	0111111111111100,
	16'b	0010000011111110,
	16'b	0000000001111110,
	16'b	0000000000111111,
	16'b	0000000000011111,
	16'b	0000000000011111,
	16'b	0000000000001111,
	16'b	0000000000001111,
	16'b	0000000000001111,
	16'b	0000000000011111,
	16'b	0000000000011111,
	16'b	1000000000111110,
	16'b	1100000001111110,
	16'b	1111100011111100,
	16'b	1111111111111000,
	16'b	1111111111111000,
	16'b	1111111111110000,
	16'b	0001111111000000},
																		
	{16'b	0000000111111100,
	16'b	0000011111111110,
	16'b	0000111111111110,
	16'b	0001111111111111,
	16'b	0001111100001111,
	16'b	0011111100000001,
	16'b	0011111000000000,
	16'b	0111110000000000,
	16'b	0111100000000000,
	16'b	1111100000000000,
	16'b	1111000000000000,
	16'b	1111000000000000,
	16'b	1111000000000000,
	16'b	1111001111111000,
	16'b	1111111111111100,
	16'b	1111111111111110,
	16'b	1111111111111111,
	16'b	1111111101111111,
	16'b	1111100000011111,
	16'b	1111000000001111,
	16'b	1111000000000111,
	16'b	1111000000000111,
	16'b	1111000000000111,
	16'b	1111000000000111,
	16'b	1111100000001111,
	16'b	1111100000001111,
	16'b	0111110000011111,
	16'b	0111111101111110,
	16'b	0011111111111110,
	16'b	0001111111111100,
	16'b	0001111111111000,
	16'b	0000011111100000},
																		
	{16'b	1111111111111111,
	16'b	1111111111111111,
	16'b	1111111111111111,
	16'b	1111111111111111,
	16'b	1100000000001111,
	16'b	1000000000011111,
	16'b	0000000000011111,
	16'b	0000000000011110,
	16'b	0000000000111110,
	16'b	0000000000111100,
	16'b	0000000001111100,
	16'b	0000000001111000,
	16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0000000011111000,
	16'b	0000000011110000,
	16'b	0000000011110000,
	16'b	0000000011100000,
	16'b	0000000011100000,
	16'b	0000000111100000,
	16'b	0000000111100000,
	16'b	0000001111000000,
	16'b	0000001111000000,
	16'b	0000011110000000,
	16'b	0000011110000000,
	16'b	0000111110000000,
	16'b	0000111100000000,
	16'b	0000111100000000,
	16'b	0001111100000000,
	16'b	0001111100000000,
	16'b	0001111100000000},
																		
	{16'b	0000111111110000,
	16'b	0001111111111000,
	16'b	0011111111111100,
	16'b	0111111111111110,
	16'b	0111111011111110,
	16'b	1111100000111111,
	16'b	1111100000011111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111000000001111,
	16'b	1111100000011110,
	16'b	0111110000111110,
	16'b	0111111001111100,
	16'b	0011111111111000,
	16'b	0001111111111000,
	16'b	0000111111100000,
	16'b	0000111111110000,
	16'b	0001111111111000,
	16'b	0011111111111100,
	16'b	0111111001111110,
	16'b	1111100000111111,
	16'b	1111000000001111,
	16'b	1110000000001111,
	16'b	1110000000000111,
	16'b	1110000000000111,
	16'b	1111000000001111,
	16'b	1111100000011111,
	16'b	1111111001111111,
	16'b	1111111111111110,
	16'b	0111111111111110,
	16'b	0011111111111000,
	16'b	0001111111110000},
																		
	{16'b	0000111111100000,
	16'b	0001111111111000,
	16'b	0011111111111000,
	16'b	0111111111111100,
	16'b	1111111011111100,
	16'b	1111100000111110,
	16'b	1111000000011110,
	16'b	1111000000011111,
	16'b	1110000000001111,
	16'b	1110000000001111,
	16'b	1110000000001111,
	16'b	1110000000001111,
	16'b	1111000000001111,
	16'b	1111100000011111,
	16'b	1111111011111111,
	16'b	1111111111111111,
	16'b	0111111111111111,
	16'b	0011111111111111,
	16'b	0001111111001111,
	16'b	0000000000001111,
	16'b	0000000000001111,
	16'b	0000000000001111,
	16'b	0000000000011110,
	16'b	0000000000011110,
	16'b	0000000000111110,
	16'b	0000000001111100,
	16'b	1000000011111100,
	16'b	1111000011111000,
	16'b	1111111111111000,
	16'b	1111111111110000,
	16'b	1111111111100000,
	16'b	0011111100000000},

};
 
// assign offsetY_LSB  = offsetY[4:0] ; // get lower 5 bits 
// assign offsetY_MSB  = offsetY[8:5] ; // get higher 4 bits 
// assign offsetX_LSB  = offsetX[4:0] ; 
// assign offsetX_MSB  = offsetX[8:5] ; 

// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBitMapMask  <=  MazeDefaultBitMapMask ;  //  copy default tabel 
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 
//----------------------------------add collision betwenn smiley and Hart -- disappear Hart  ------------------------------------------		
             if (smiley_hart_collision == 1'b1)
						MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h0;


		
//------------------------------------End collision betwenn smiley and Hart-------------------------------------------- 		
		
		if (InsideRectangle == 1'b1 )	
			begin 
		   	case (MazeBitMapMask[offsetY[8:5]][offsetX[8:5]])
					 4'h0 : RGBout <= TRANSPARENT_ENCODING ;
					 4'h1 : RGBout <= object_colors[random_hart][offsetY[4:0]][offsetX[4:0]]; 
					 4'h2 : RGBout <= object_colors[2'h1][offsetY[4:0]][offsetX[4:0]] ; 
					 default:  RGBout <= TRANSPARENT_ENCODING ; 
				endcase
			end 
 
	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

